----------------------------------------------------------------------------------
-- COMPANY: 
-- ENGINEER: 
-- 
-- CREATE DATE:    17:03:25 11/13/2019 
-- DESIGN NAME: 
-- MODULE NAME:    BCD_CHECKER - BEHAVIORAL 
-- PROJECT NAME: 
-- TARGET DEVICES: 
-- TOOL VERSIONS: 
-- DESCRIPTION: 
--
-- DEPENDENCIES: 
--
-- REVISION: 
-- REVISION 0.01 - FILE CREATED
-- ADDITIONAL COMMENTS: 
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF USING
-- ARITHMETIC FUNCTIONS WITH SIGNED OR UNSIGNED VALUES
--USE IEEE.NUMERIC_STD.ALL;

-- UNCOMMENT THE FOLLOWING LIBRARY DECLARATION IF INSTANTIATING
-- ANY XILINX PRIMITIVES IN THIS CODE.
--LIBRARY UNISIM;
--USE UNISIM.VCOMPONENTS.ALL;

ENTITY CHECK_BCD IS
PORT(

N1: IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
N2: IN STD_LOGIC_VECTOR (3 DOWNTO 0);

K: OUT STD_LOGIC



);
END CHECK_BCD;

ARCHITECTURE BEHAVIORAL OF CHECK_BCD IS

BEGIN

PROCESS(N1, N2)

BEGIN

IF(N1>"1001" OR N2>"1001" OR  (N2="0000" AND N1="0000")) THEN 
	K<='0';
ELSE  
	K<='1';
END IF ;


END PROCESS;



END BEHAVIORAL;

